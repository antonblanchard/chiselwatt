module Chiselwatt_pll(
  input  clki,
  output clko,
  output lock
);
  (* ICP_CURRENT="12" *) (* LPF_RESISTOR="8" *) (* MFG_ENABLE_FILTEROPAMP="1" *) (* MFG_GMCREF_SEL="2" *)

  EHXPLLL #(
    .PLLRST_ENA("DISABLED"),
    .INTFB_WAKE("DISABLED"),
    .STDBY_ENABLE("DISABLED"),
    .DPHASE_SOURCE("DISABLED"),
    .CLKOP_FPHASE(0),
    .CLKOP_CPHASE(11),
    .OUTDIVIDER_MUXA("DIVA"),
    .CLKOP_ENABLE("ENABLED"),
    .CLKOP_DIV(12),
    .CLKFB_DIV(25),
    .CLKI_DIV(6),
    .FEEDBK_PATH("CLKOP")
  ) pll_i (
    .CLKI(clki),
    .CLKFB(clko),
    .CLKOP(clko),
    .LOCK(lock),
    .RST(1'b0),
    .STDBY(1'b0),
    .PHASESEL0(1'b0),
    .PHASESEL1(1'b0),
    .PHASEDIR(1'b0),
    .PHASESTEP(1'b0),
    .PLLWAKESYNC(1'b0),
    .ENCLKOP(1'b0)
  );

endmodule
